`timescale 1ns / 1ps

module Mux4Way16_tb();

    reg [15:0] a;
    reg [15:0] b;
    reg [15:0] c;
    reg [15:0] d;
    reg [1:0] sel;
    wire [15:0] out;

    Mux4Way16 u_Mux4Way16(
        .a_i(a),
        .b_i(b),
        .c_i(c),
        .d_i(d),
        .sel_i(sel),
        .out_o(out)
    );

    initial begin
        a = 16'b0000_0000_0000_0000;b = 16'b0000_0000_0000_0000;
        c = 16'b0000_0000_0000_0000;d = 16'b0000_0000_0000_0000;
        sel = 2'b00;
        $display("test running...");
        #10
        a = 16'b0000_0000_0000_0000;b = 16'b0000_0000_0000_0000;
        c = 16'b0000_0000_0000_0000;d = 16'b0000_0000_0000_0000;
        sel = 2'b00;
        #10
        a = 16'b0000_0000_0000_0000;b = 16'b0000_0000_0000_0000;
        c = 16'b0000_0000_0000_0000;d = 16'b0000_0000_0000_0000;
        sel = 2'b01;
        #10
        a = 16'b0000_0000_0000_0000;b = 16'b0000_0000_0000_0000;
        c = 16'b0000_0000_0000_0000;d = 16'b0000_0000_0000_0000;
        sel = 2'b10;
        #10
        a = 16'b0000_0000_0000_0000;b = 16'b0000_0000_0000_0000;
        c = 16'b0000_0000_0000_0000;d = 16'b0000_0000_0000_0000;
        sel = 2'b11;
        #10
        a = 16'b0001001000110100;b = 16'b1001100001110110;
        c = 16'b1010101010101010;d = 16'b0101010101010101;
        sel = 2'b00;
        #10
        a = 16'b0001001000110100;b = 16'b1001100001110110;
        c = 16'b1010101010101010;d = 16'b0101010101010101;
        sel = 2'b01;
        #10
        a = 16'b0001001000110100;b = 16'b1001100001110110;
        c = 16'b1010101010101010;d = 16'b0101010101010101;
        sel = 2'b10;
        #10
        a = 16'b0001001000110100;b = 16'b1001100001110110;
        c = 16'b1010101010101010;d = 16'b0101010101010101;
        sel = 2'b11;
        #1000 
        $finish;
    end

    initial begin
        $dumpfile("vtest/dumpfile/Mux4Way16.vcd");
	    $dumpvars(0,Mux4Way16_tb);
	end

endmodule