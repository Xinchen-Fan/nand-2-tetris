`timescale 1ns / 1ps

module Mux8Way16_tb();

    reg [15:0] a;
    reg [15:0] b;
    reg [15:0] c;
    reg [15:0] d;
    reg [15:0] e;
    reg [15:0] f;
    reg [15:0] g;
    reg [15:0] h;
    reg [2:0] sel;
    wire [15:0] out;

    Mux8Way16 u_Mux8Way16(
        .a_i(a),
        .b_i(b),
        .c_i(c),
        .d_i(d),
        .e_i(e),
        .f_i(f),
        .g_i(g),
        .h_i(h),
        .sel_i(sel),
        .out_o(out)
    );

    initial begin
        a = 16'b0000_0000_0000_0000;b = 16'b0000_0000_0000_0000;
        c = 16'b0000_0000_0000_0000;d = 16'b0000_0000_0000_0000;
        e = 16'b0000_0000_0000_0000;f = 16'b0000_0000_0000_0000;
        g = 16'b0000_0000_0000_0000;h = 16'b0000_0000_0000_0000;
        sel = 3'b000;
        $display("test running...");
        #10
        a = 16'b0000_0000_0000_0000;b = 16'b0000_0000_0000_0000;
        c = 16'b0000_0000_0000_0000;d = 16'b0000_0000_0000_0000;
        e = 16'b0000_0000_0000_0000;f = 16'b0000_0000_0000_0000;
        g = 16'b0000_0000_0000_0000;h = 16'b0000_0000_0000_0000;
        sel = 3'b000;
        #10 sel = 3'b001;
        #10 sel = 3'b010;
        #10 sel = 3'b011;
        #10 sel = 3'b100;
        #10 sel = 3'b101;
        #10 sel = 3'b110;
        #10 sel = 3'b111;
        #10
        a = 16'b0001001000110100;b = 16'b0010001101000101;
        c = 16'b0011010001010110;d = 16'b0100010101100111;
        e = 16'b0101011001111000;f = 16'b0110011110001001;
        g = 16'b0111100010011010;h = 16'b1000100110101011;
        sel = 3'b000;
        #10 sel = 3'b001;
        #10 sel = 3'b010;
        #10 sel = 3'b011;
        #10 sel = 3'b100;
        #10 sel = 3'b101;
        #10 sel = 3'b110;
        #10 sel = 3'b111;
        #1000 
        $finish;
    end

    initial begin
        $dumpfile("vtest/dumpfile/Mux8Way16.vcd");
	    $dumpvars(0,Mux8Way16_tb);
	end

endmodule