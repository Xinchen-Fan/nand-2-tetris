/* Program Counter

 * A 16-bit counter with load and reset control bits.
 * if      (reset[t] == 1) out[t+1] = 0
 * else if (load[t] == 1)  out[t+1] = in[t]
 * else if (inc[t] == 1)   out[t+1] = out[t] + 1  (integer addition)
 * else                    out[t+1] = out[t]

PC u_PC(
    .clk_i(),
    .in_i(),
    .load_i(),
    .inc_i(),
    .reset_i(),
    .out_o()
);


 */

 module PC(
    input wire clk_i,
    input wire [15:0] in_i,
    input wire load_i,
    input wire inc_i,
    input wire reset_i,
    output wire [15:0] out_o
);

    wire [15:0] in_inc;
    wire [15:0] in_tmp1;
    wire [15:0] in_tmp2;
    wire [15:0] in_new;
    wire [15:0] out_buf;
    assign out_o = out_buf;

    assign in_inc = out_buf + 1'b1; // pc+1
    assign in_tmp1 = inc_i ? in_inc : out_buf; // +1 or hold
    assign in_tmp2 = load_i ? in_i : in_tmp1;  // load or (+1 or hold)
    // assign in_new = reset_i ? 16'b0 : in_tmp2; // reset or (load or (+1 or hold))

    Register #(16, 16'b0) u_Register(.clk_i(clk_i), .in_i(in_tmp2), .reset_i(reset_i), .load_i(1'b1), .out_o(out_buf));


endmodule

